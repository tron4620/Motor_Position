
module sysPll (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
